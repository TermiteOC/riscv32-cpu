-------------------------------------------------------------------------------
-- Module: ALU_1Bit
-- Description:
--   - 1-bit ALU supporting AND, OR, ADD, SUB, NOR, NAND operations.
--   - Supports SLT operation only if it is paired with other 1-bit ALUs
--   - Supports input inversion for a and b to enable complementary operations.
-- Author: Levy Elmescany
-- Date: 2025-07-24
-- License: MIT
-- Inputs: a, b, cin, less, a_invert, b_invert, op
-- Outputs: res, cout
-- Tool Compatibility: Quartus Prime 24.x or compatible synthesis tools
-- Notes:
--   - Uses internal components:
--     - 2-to-1 multiplexer for selecting NOT a or NOT b
--     - 4-to-1 multiplexer for operation
--     - Full adder
--   - a_invert and b_invert control input inversion.
--   - NAND and NOR are generated by inverting inputs and using OR/AND operations.
--   - Less input and set output are only used in the SLT operation:
--     - Set is computed in MSB and indicates a < b result
--     - Less is used in LSB to select res = set
-- Simulation: None (to be tested via ALU_32Bit simulation)
-- Revision History:
--   Rev 1.0 - 2025-07-24 - Initial implementation
--   Rev 1.1 - 2025-07-27 - Syntax fix: removed extra semicolon in entity port declaration
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ALU_1Bit is
    port (
        a        : in  std_logic;                    -- 1st operand
        b        : in  std_logic;                    -- 2nd operand
        cin      : in  std_logic;                    -- carry-in
        less     : in  std_logic;                    -- value if a is less than b (LSB)
        a_invert : in  std_logic;                    -- inverted a selector
        b_invert : in  std_logic;                    -- inverted b selector
        op       : in  std_logic_vector(1 downto 0); -- operation selector
        res      : out std_logic;                    -- result
        cout     : out std_logic;                    -- carry-out from adder
        set      : out std_logic                     -- sets value if a is less than b (MSB)
    );
end ALU_1Bit;

architecture rtl of ALU_1Bit is

    -- 1-bit 2-to-1 multiplexer
    component Mux2x1_1Bit is
        port (
            sel    : in  std_logic;                    -- selector
            inputs : in  std_logic_vector(1 downto 0); -- 2 inputs
            output : out std_logic;                    -- 1 output
        );
    end component;

    -- 1-bit full adder
    component FullAdder_1Bit is
        port (
            a    : in  std_logic; -- 1st operand
            b    : in  std_logic; -- 2nd operand
            cin  : in  std_logic; -- carry-in
            sum  : out std_logic; -- result of the sum
            cout : out std_logic  -- carry-out
        );
    end component;

    -- 1-bit 4-to-1 multiplexer
    component Mux4x1_1Bit is
        port (
            sel    : in  std_logic_vector(1 downto 0); -- selector
            inputs : in  std_logic_vector(3 downto 0); -- 4 inputs
            output : out std_logic;                    -- 1 output
        );
    end component;
    
    -- Vector input for inverted muxes
    signal w_a_mux_in : std_logic_vector(1 downto 0);
    signal w_b_mux_in : std_logic_vector(1 downto 0);
    
    -- Output of the inverted muxes
    signal w_a_mux_out : std_logic;
    signal w_b_mux_out : std_logic;

    -- Operation results
    signal w_and : std_logic;
    signal w_or  : std_logic;
    signal w_sum : std_logic;
    
    -- Carry-out from the adder
    signal w_cout : std_logic;

    -- Overflow detector signal
    signal w_overflow : std_logic;

    -- Vector input for the 4-to-1 mux
    signal w_op_mux_in : std_logic_vector(3 downto 0);

begin
    -- Combinational Logic
    -- Input vectors for muxes: bit 0 = original input, bit 1 = inverted input
    w_a_mux_in(0) <= a;
    w_a_mux_in(1) <= not a;
    w_b_mux_in(0) <= b;
    w_b_mux_in(1) <= not b;

    w_and <= w_a_mux_out and w_b_mux_out;
    w_or  <= w_a_mux_out or w_b_mux_out;

    -- If the carry-in and carry-out of MSB is different, overflow exists
    w_overflow <= cin xor w_cout;

    -- Set is 1 if the sign of the sum is negative, but if overflow is 1, the sign inverts
    set <= w_sum xor w_overflow;

    -- Mux inputs indexed as: 0 = AND, 1 = OR, 2 = SUM, 3 = SLT
    w_op_mux_in(0) <= w_and;
    w_op_mux_in(1) <= w_or;
    w_op_mux_in(2) <= w_sum;
    w_op_mux_in(3) <= less;

    -- Component Instantiations
    -- Multiplexer that selects original a or inverted a. Selector: 0 = original, 1 = inverted
    mux2x1_a_inst : Mux2x1_1Bit
    port map (
        sel    => a_invert,
        inputs => w_a_mux_in,
        output => w_a_mux_out
    );

    -- Multiplexer that selects original b or inverted b. Selector: 0 = original, 1 = inverted
    mux2x1_b_inst : Mux2x1_1Bit
    port map (
        sel    => b_invert,
        inputs => w_b_mux_in,
        output => w_b_mux_out
    );

    full_adder_inst : FullAdder_1Bit 
    port map (
        a    => w_a_mux_out,
        b    => w_b_mux_out,
        cin  => cin,
        sum  => w_sum,
        cout => w_cout
    );
    
    -- Multiplexer that selects operation. Selector: 00 = AND, 01 = OR, 10 = ADD, 11 = SLT
    mux4x1_inst : Mux4x1_1Bit
    port map (
        sel    => op,
        inputs => w_op_mux_in,
        output => res
    );
end rtl;