library IEEE;
use IEEE.std_logic_1164.all;

package CommonTypes is
    -- Shared types
    type WordArray_t is array(0 to 31) of std_logic_vector(31 downto 0);
end package;

package body CommonTypes is
end package body;
